package exec_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "exec_seq_item.svh"
typedef uvm_sequencer #(exec_seq_item) exec_sequencer;
`include "exec_agent_config.svh"
`include "exec_driver.svh"
//`include "exec_coverage_monitor.svh"
`include "exec_monitor.svh"
`include "exec_agent.svh"

// Utility Sequences
`include "exec_seq.svh"

endpackage
