// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package cosim_agent_pkg;
  import uvm_pkg::*;


  `include "uvm_macros.svh"
  `include "spike_cosim_dpi.svh"
  `include "cosim_dpi.svh"
  
endpackage
