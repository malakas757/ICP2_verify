package fetch_env_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import bpu_agent_pkg::*;
	import exec_agent_pkg::*;
	import if_id_agent_pkg::*;
	
	`include "fetch_env_config.svh"
	`include "refmod.svh"
	`include "if_scoreboard.svh"
	`include "fetch_env.svh"




endpackage
