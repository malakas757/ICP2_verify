package if_id_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "if_id_seq_item.svh"
//typedef uvm_sequencer #(if_id_seq_item) if_id_sequencer;
`include "if_id_agent_config.svh"
//`include "if_id_driver.svh"
//`include "if_id_coverage_monitor.svh"
`include "if_id_monitor.svh"
`include "if_id_agent.svh"

// Utility Sequences
//`include "if_id_seq.svh"

endpackage
