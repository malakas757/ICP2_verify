package fetch_vseq_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	import bpu_agent_pkg::*;
	import exec_agent_pkg::*;
	import seq_pkg::*;

	
	`include "fetch_vseq_base.svh"
	`include "fetch_random_vseq.svh"
endpackage