interface bpu_if(input clk, input rstn);
    logic pred;

endinterface